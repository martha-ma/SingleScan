// kernel.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module kernel (
		input  wire [3:0]  alarm_select_export,     //      alarm_select.export
		input  wire        clk_clk,                 //               clk.clk
		output wire        epcs_flash_dclk,         //        epcs_flash.dclk
		output wire        epcs_flash_sce,          //                  .sce
		output wire        epcs_flash_sdo,          //                  .sdo
		input  wire        epcs_flash_data0,        //                  .data0
		input  wire        laser_fifo_in_valid,     //     laser_fifo_in.valid
		input  wire [31:0] laser_fifo_in_data,      //                  .data
		output wire        laser_fifo_in_ready,     //                  .ready
		output wire        power_led_export,        //         power_led.export
		output wire        protocol_fifo_out_valid, // protocol_fifo_out.valid
		output wire [31:0] protocol_fifo_out_data,  //                  .data
		input  wire        protocol_fifo_out_ready, //                  .ready
		input  wire        reset_reset_n,           //             reset.reset_n
		output wire        scl_export,              //               scl.export
		inout  wire        sda_export,              //               sda.export
		input  wire        spird_fifo_in_valid,     //     spird_fifo_in.valid
		input  wire [31:0] spird_fifo_in_data,      //                  .data
		output wire        spird_fifo_in_ready,     //                  .ready
		output wire        spiwr_fifo_out_valid,    //    spiwr_fifo_out.valid
		output wire [31:0] spiwr_fifo_out_data,     //                  .data
		input  wire        spiwr_fifo_out_ready,    //                  .ready
		output wire        status_led_export,       //        status_led.export
		output wire        w5500_cs_export,         //          w5500_cs.export
		input  wire        w5500_int_in_port,       //         w5500_int.in_port
		output wire        w5500_int_out_port,      //                  .out_port
		output wire        w5500_rst_export         //         w5500_rst.export
	);

	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                             // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [19:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [19:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                    // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;          // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;       // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;           // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;              // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;             // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_epcs_control_port_chipselect -> epcs_flash:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_readdata;   // epcs_flash:readdata -> mm_interconnect_0:epcs_flash_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_epcs_control_port_address -> epcs_flash:address
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_epcs_control_port_read -> epcs_flash:read_n
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_epcs_control_port_write -> epcs_flash:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_epcs_control_port_writedata -> epcs_flash:writedata
	wire         mm_interconnect_0_protocol_fifo_in_waitrequest;            // protocol_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_0:protocol_fifo_in_waitrequest
	wire   [0:0] mm_interconnect_0_protocol_fifo_in_address;                // mm_interconnect_0:protocol_fifo_in_address -> protocol_fifo:avalonmm_write_slave_address
	wire         mm_interconnect_0_protocol_fifo_in_write;                  // mm_interconnect_0:protocol_fifo_in_write -> protocol_fifo:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_protocol_fifo_in_writedata;              // mm_interconnect_0:protocol_fifo_in_writedata -> protocol_fifo:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_spiwr_fifo_in_waitrequest;               // spiwr_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_0:spiwr_fifo_in_waitrequest
	wire   [0:0] mm_interconnect_0_spiwr_fifo_in_address;                   // mm_interconnect_0:spiwr_fifo_in_address -> spiwr_fifo:avalonmm_write_slave_address
	wire         mm_interconnect_0_spiwr_fifo_in_write;                     // mm_interconnect_0:spiwr_fifo_in_write -> spiwr_fifo:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_spiwr_fifo_in_writedata;                 // mm_interconnect_0:spiwr_fifo_in_writedata -> spiwr_fifo:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_laser_fifo_in_csr_readdata;              // laser_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:laser_fifo_in_csr_readdata
	wire   [2:0] mm_interconnect_0_laser_fifo_in_csr_address;               // mm_interconnect_0:laser_fifo_in_csr_address -> laser_fifo:wrclk_control_slave_address
	wire         mm_interconnect_0_laser_fifo_in_csr_read;                  // mm_interconnect_0:laser_fifo_in_csr_read -> laser_fifo:wrclk_control_slave_read
	wire         mm_interconnect_0_laser_fifo_in_csr_write;                 // mm_interconnect_0:laser_fifo_in_csr_write -> laser_fifo:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_laser_fifo_in_csr_writedata;             // mm_interconnect_0:laser_fifo_in_csr_writedata -> laser_fifo:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_protocol_fifo_in_csr_readdata;           // protocol_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:protocol_fifo_in_csr_readdata
	wire   [2:0] mm_interconnect_0_protocol_fifo_in_csr_address;            // mm_interconnect_0:protocol_fifo_in_csr_address -> protocol_fifo:wrclk_control_slave_address
	wire         mm_interconnect_0_protocol_fifo_in_csr_read;               // mm_interconnect_0:protocol_fifo_in_csr_read -> protocol_fifo:wrclk_control_slave_read
	wire         mm_interconnect_0_protocol_fifo_in_csr_write;              // mm_interconnect_0:protocol_fifo_in_csr_write -> protocol_fifo:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_protocol_fifo_in_csr_writedata;          // mm_interconnect_0:protocol_fifo_in_csr_writedata -> protocol_fifo:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_spiwr_fifo_in_csr_readdata;              // spiwr_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:spiwr_fifo_in_csr_readdata
	wire   [2:0] mm_interconnect_0_spiwr_fifo_in_csr_address;               // mm_interconnect_0:spiwr_fifo_in_csr_address -> spiwr_fifo:wrclk_control_slave_address
	wire         mm_interconnect_0_spiwr_fifo_in_csr_read;                  // mm_interconnect_0:spiwr_fifo_in_csr_read -> spiwr_fifo:wrclk_control_slave_read
	wire         mm_interconnect_0_spiwr_fifo_in_csr_write;                 // mm_interconnect_0:spiwr_fifo_in_csr_write -> spiwr_fifo:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_spiwr_fifo_in_csr_writedata;             // mm_interconnect_0:spiwr_fifo_in_csr_writedata -> spiwr_fifo:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_spird_fifo_in_csr_readdata;              // spird_fifo:wrclk_control_slave_readdata -> mm_interconnect_0:spird_fifo_in_csr_readdata
	wire   [2:0] mm_interconnect_0_spird_fifo_in_csr_address;               // mm_interconnect_0:spird_fifo_in_csr_address -> spird_fifo:wrclk_control_slave_address
	wire         mm_interconnect_0_spird_fifo_in_csr_read;                  // mm_interconnect_0:spird_fifo_in_csr_read -> spird_fifo:wrclk_control_slave_read
	wire         mm_interconnect_0_spird_fifo_in_csr_write;                 // mm_interconnect_0:spird_fifo_in_csr_write -> spird_fifo:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_spird_fifo_in_csr_writedata;             // mm_interconnect_0:spird_fifo_in_csr_writedata -> spird_fifo:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_spird_fifo_out_readdata;                 // spird_fifo:avalonmm_read_slave_readdata -> mm_interconnect_0:spird_fifo_out_readdata
	wire         mm_interconnect_0_spird_fifo_out_waitrequest;              // spird_fifo:avalonmm_read_slave_waitrequest -> mm_interconnect_0:spird_fifo_out_waitrequest
	wire   [0:0] mm_interconnect_0_spird_fifo_out_address;                  // mm_interconnect_0:spird_fifo_out_address -> spird_fifo:avalonmm_read_slave_address
	wire         mm_interconnect_0_spird_fifo_out_read;                     // mm_interconnect_0:spird_fifo_out_read -> spird_fifo:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_laser_fifo_out_readdata;                 // laser_fifo:avalonmm_read_slave_readdata -> mm_interconnect_0:laser_fifo_out_readdata
	wire         mm_interconnect_0_laser_fifo_out_waitrequest;              // laser_fifo:avalonmm_read_slave_waitrequest -> mm_interconnect_0:laser_fifo_out_waitrequest
	wire   [0:0] mm_interconnect_0_laser_fifo_out_address;                  // mm_interconnect_0:laser_fifo_out_address -> laser_fifo:avalonmm_read_slave_address
	wire         mm_interconnect_0_laser_fifo_out_read;                     // mm_interconnect_0:laser_fifo_out_read -> laser_fifo:avalonmm_read_slave_read
	wire         mm_interconnect_0_w5500_rst_s1_chipselect;                 // mm_interconnect_0:w5500_rst_s1_chipselect -> w5500_rst:chipselect
	wire  [31:0] mm_interconnect_0_w5500_rst_s1_readdata;                   // w5500_rst:readdata -> mm_interconnect_0:w5500_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_w5500_rst_s1_address;                    // mm_interconnect_0:w5500_rst_s1_address -> w5500_rst:address
	wire         mm_interconnect_0_w5500_rst_s1_write;                      // mm_interconnect_0:w5500_rst_s1_write -> w5500_rst:write_n
	wire  [31:0] mm_interconnect_0_w5500_rst_s1_writedata;                  // mm_interconnect_0:w5500_rst_s1_writedata -> w5500_rst:writedata
	wire         mm_interconnect_0_w5500_int_s1_chipselect;                 // mm_interconnect_0:w5500_int_s1_chipselect -> w5500_int:chipselect
	wire  [31:0] mm_interconnect_0_w5500_int_s1_readdata;                   // w5500_int:readdata -> mm_interconnect_0:w5500_int_s1_readdata
	wire   [1:0] mm_interconnect_0_w5500_int_s1_address;                    // mm_interconnect_0:w5500_int_s1_address -> w5500_int:address
	wire         mm_interconnect_0_w5500_int_s1_write;                      // mm_interconnect_0:w5500_int_s1_write -> w5500_int:write_n
	wire  [31:0] mm_interconnect_0_w5500_int_s1_writedata;                  // mm_interconnect_0:w5500_int_s1_writedata -> w5500_int:writedata
	wire         mm_interconnect_0_w5500_cs_s1_chipselect;                  // mm_interconnect_0:w5500_cs_s1_chipselect -> w5500_cs:chipselect
	wire  [31:0] mm_interconnect_0_w5500_cs_s1_readdata;                    // w5500_cs:readdata -> mm_interconnect_0:w5500_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_w5500_cs_s1_address;                     // mm_interconnect_0:w5500_cs_s1_address -> w5500_cs:address
	wire         mm_interconnect_0_w5500_cs_s1_write;                       // mm_interconnect_0:w5500_cs_s1_write -> w5500_cs:write_n
	wire  [31:0] mm_interconnect_0_w5500_cs_s1_writedata;                   // mm_interconnect_0:w5500_cs_s1_writedata -> w5500_cs:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_scl_s1_chipselect;                       // mm_interconnect_0:SCL_s1_chipselect -> SCL:chipselect
	wire  [31:0] mm_interconnect_0_scl_s1_readdata;                         // SCL:readdata -> mm_interconnect_0:SCL_s1_readdata
	wire   [1:0] mm_interconnect_0_scl_s1_address;                          // mm_interconnect_0:SCL_s1_address -> SCL:address
	wire         mm_interconnect_0_scl_s1_write;                            // mm_interconnect_0:SCL_s1_write -> SCL:write_n
	wire  [31:0] mm_interconnect_0_scl_s1_writedata;                        // mm_interconnect_0:SCL_s1_writedata -> SCL:writedata
	wire         mm_interconnect_0_sda_s1_chipselect;                       // mm_interconnect_0:SDA_s1_chipselect -> SDA:chipselect
	wire  [31:0] mm_interconnect_0_sda_s1_readdata;                         // SDA:readdata -> mm_interconnect_0:SDA_s1_readdata
	wire   [1:0] mm_interconnect_0_sda_s1_address;                          // mm_interconnect_0:SDA_s1_address -> SDA:address
	wire         mm_interconnect_0_sda_s1_write;                            // mm_interconnect_0:SDA_s1_write -> SDA:write_n
	wire  [31:0] mm_interconnect_0_sda_s1_writedata;                        // mm_interconnect_0:SDA_s1_writedata -> SDA:writedata
	wire         mm_interconnect_0_power_led_s1_chipselect;                 // mm_interconnect_0:power_led_s1_chipselect -> power_led:chipselect
	wire  [31:0] mm_interconnect_0_power_led_s1_readdata;                   // power_led:readdata -> mm_interconnect_0:power_led_s1_readdata
	wire   [1:0] mm_interconnect_0_power_led_s1_address;                    // mm_interconnect_0:power_led_s1_address -> power_led:address
	wire         mm_interconnect_0_power_led_s1_write;                      // mm_interconnect_0:power_led_s1_write -> power_led:write_n
	wire  [31:0] mm_interconnect_0_power_led_s1_writedata;                  // mm_interconnect_0:power_led_s1_writedata -> power_led:writedata
	wire         mm_interconnect_0_status_led_s1_chipselect;                // mm_interconnect_0:status_led_s1_chipselect -> status_led:chipselect
	wire  [31:0] mm_interconnect_0_status_led_s1_readdata;                  // status_led:readdata -> mm_interconnect_0:status_led_s1_readdata
	wire   [1:0] mm_interconnect_0_status_led_s1_address;                   // mm_interconnect_0:status_led_s1_address -> status_led:address
	wire         mm_interconnect_0_status_led_s1_write;                     // mm_interconnect_0:status_led_s1_write -> status_led:write_n
	wire  [31:0] mm_interconnect_0_status_led_s1_writedata;                 // mm_interconnect_0:status_led_s1_writedata -> status_led:writedata
	wire         mm_interconnect_0_led_timer_s1_chipselect;                 // mm_interconnect_0:led_timer_s1_chipselect -> led_timer:chipselect
	wire  [15:0] mm_interconnect_0_led_timer_s1_readdata;                   // led_timer:readdata -> mm_interconnect_0:led_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_led_timer_s1_address;                    // mm_interconnect_0:led_timer_s1_address -> led_timer:address
	wire         mm_interconnect_0_led_timer_s1_write;                      // mm_interconnect_0:led_timer_s1_write -> led_timer:write_n
	wire  [15:0] mm_interconnect_0_led_timer_s1_writedata;                  // mm_interconnect_0:led_timer_s1_writedata -> led_timer:writedata
	wire         mm_interconnect_0_alarm_select_s1_chipselect;              // mm_interconnect_0:alarm_select_s1_chipselect -> alarm_select:chipselect
	wire  [31:0] mm_interconnect_0_alarm_select_s1_readdata;                // alarm_select:readdata -> mm_interconnect_0:alarm_select_s1_readdata
	wire   [1:0] mm_interconnect_0_alarm_select_s1_address;                 // mm_interconnect_0:alarm_select_s1_address -> alarm_select:address
	wire         mm_interconnect_0_alarm_select_s1_write;                   // mm_interconnect_0:alarm_select_s1_write -> alarm_select:write_n
	wire  [31:0] mm_interconnect_0_alarm_select_s1_writedata;               // mm_interconnect_0:alarm_select_s1_writedata -> alarm_select:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // epcs_flash:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // led_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // alarm_select:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_irq_irq;                                             // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [SCL:reset_n, SDA:reset_n, alarm_select:reset_n, epcs_flash:reset_n, irq_mapper:reset, jtag_uart:rst_n, led_timer:reset_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, onchip_memory:reset, power_led:reset_n, protocol_fifo:reset_n, rst_translator:in_reset, spird_fifo:reset_n, spiwr_fifo:reset_n, status_led:reset_n, sysid:reset_n, w5500_cs:reset_n, w5500_int:reset_n, w5500_rst:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [epcs_flash:reset_req, nios2:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                           // nios2:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [laser_fifo:reset_n, mm_interconnect_0:laser_fifo_reset_in_reset_bridge_in_reset_reset]

	kernel_SCL scl (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scl_s1_readdata),   //                    .readdata
		.out_port   (scl_export)                           // external_connection.export
	);

	kernel_SDA sda (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sda_s1_readdata),   //                    .readdata
		.bidir_port (sda_export)                           // external_connection.export
	);

	kernel_alarm_select alarm_select (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_alarm_select_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_alarm_select_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_alarm_select_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_alarm_select_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_alarm_select_s1_readdata),   //                    .readdata
		.in_port    (alarm_select_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                      //                 irq.irq
	);

	kernel_epcs_flash epcs_flash (
		.clk        (clk_clk),                                                   //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                        //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver1_irq),                                  //               irq.irq
		.dclk       (epcs_flash_dclk),                                           //          external.export
		.sce        (epcs_flash_sce),                                            //                  .export
		.sdo        (epcs_flash_sdo),                                            //                  .export
		.data0      (epcs_flash_data0)                                           //                  .export
	);

	kernel_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	kernel_laser_fifo laser_fifo (
		.wrclock                         (clk_clk),                                       //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),           // reset_in.reset_n
		.avalonst_sink_valid             (laser_fifo_in_valid),                           //       in.valid
		.avalonst_sink_data              (laser_fifo_in_data),                            //         .data
		.avalonst_sink_ready             (laser_fifo_in_ready),                           //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_laser_fifo_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_laser_fifo_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_laser_fifo_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_laser_fifo_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_0_laser_fifo_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_0_laser_fifo_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_0_laser_fifo_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_0_laser_fifo_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_0_laser_fifo_in_csr_readdata)   //         .readdata
	);

	kernel_led_timer led_timer (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_led_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_led_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_led_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_led_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_led_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                   //   irq.irq
	);

	kernel_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	kernel_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	kernel_SCL power_led (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_power_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_power_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_power_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_power_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_power_led_s1_readdata),   //                    .readdata
		.out_port   (power_led_export)                           // external_connection.export
	);

	kernel_protocol_fifo protocol_fifo (
		.wrclock                          (clk_clk),                                          //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),                  // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_protocol_fifo_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_protocol_fifo_in_write),         //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_protocol_fifo_in_address),       //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_protocol_fifo_in_waitrequest),   //         .waitrequest
		.avalonst_source_valid            (protocol_fifo_out_valid),                          //      out.valid
		.avalonst_source_data             (protocol_fifo_out_data),                           //         .data
		.avalonst_source_ready            (protocol_fifo_out_ready),                          //         .ready
		.wrclk_control_slave_address      (mm_interconnect_0_protocol_fifo_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_protocol_fifo_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_protocol_fifo_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_protocol_fifo_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_protocol_fifo_in_csr_readdata)   //         .readdata
	);

	kernel_spird_fifo spird_fifo (
		.wrclock                         (clk_clk),                                       //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonst_sink_valid             (spird_fifo_in_valid),                           //       in.valid
		.avalonst_sink_data              (spird_fifo_in_data),                            //         .data
		.avalonst_sink_ready             (spird_fifo_in_ready),                           //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_spird_fifo_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_spird_fifo_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_spird_fifo_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_spird_fifo_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_0_spird_fifo_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_0_spird_fifo_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_0_spird_fifo_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_0_spird_fifo_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_0_spird_fifo_in_csr_readdata)   //         .readdata
	);

	kernel_spiwr_fifo spiwr_fifo (
		.wrclock                          (clk_clk),                                       //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),               // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_spiwr_fifo_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_spiwr_fifo_in_write),         //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_spiwr_fifo_in_address),       //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_spiwr_fifo_in_waitrequest),   //         .waitrequest
		.avalonst_source_valid            (spiwr_fifo_out_valid),                          //      out.valid
		.avalonst_source_data             (spiwr_fifo_out_data),                           //         .data
		.avalonst_source_ready            (spiwr_fifo_out_ready),                          //         .ready
		.wrclk_control_slave_address      (mm_interconnect_0_spiwr_fifo_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_spiwr_fifo_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_spiwr_fifo_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_spiwr_fifo_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_spiwr_fifo_in_csr_readdata)   //         .readdata
	);

	kernel_SCL status_led (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_status_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_status_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_status_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_status_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_status_led_s1_readdata),   //                    .readdata
		.out_port   (status_led_export)                           // external_connection.export
	);

	kernel_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	kernel_SCL w5500_cs (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_w5500_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_w5500_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_w5500_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_w5500_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_w5500_cs_s1_readdata),   //                    .readdata
		.out_port   (w5500_cs_export)                           // external_connection.export
	);

	kernel_w5500_int w5500_int (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_w5500_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_w5500_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_w5500_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_w5500_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_w5500_int_s1_readdata),   //                    .readdata
		.in_port    (w5500_int_in_port),                         // external_connection.export
		.out_port   (w5500_int_out_port)                         //                    .export
	);

	kernel_SCL w5500_rst (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_w5500_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_w5500_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_w5500_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_w5500_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_w5500_rst_s1_readdata),   //                    .readdata
		.out_port   (w5500_rst_export)                           // external_connection.export
	);

	kernel_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                     (clk_clk),                                                   //                                   clk_clk.clk
		.laser_fifo_reset_in_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // laser_fifo_reset_in_reset_bridge_in_reset.reset
		.nios2_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                            //         nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                       (nios2_data_master_address),                                 //                         nios2_data_master.address
		.nios2_data_master_waitrequest                   (nios2_data_master_waitrequest),                             //                                          .waitrequest
		.nios2_data_master_byteenable                    (nios2_data_master_byteenable),                              //                                          .byteenable
		.nios2_data_master_read                          (nios2_data_master_read),                                    //                                          .read
		.nios2_data_master_readdata                      (nios2_data_master_readdata),                                //                                          .readdata
		.nios2_data_master_write                         (nios2_data_master_write),                                   //                                          .write
		.nios2_data_master_writedata                     (nios2_data_master_writedata),                               //                                          .writedata
		.nios2_data_master_debugaccess                   (nios2_data_master_debugaccess),                             //                                          .debugaccess
		.nios2_instruction_master_address                (nios2_instruction_master_address),                          //                  nios2_instruction_master.address
		.nios2_instruction_master_waitrequest            (nios2_instruction_master_waitrequest),                      //                                          .waitrequest
		.nios2_instruction_master_read                   (nios2_instruction_master_read),                             //                                          .read
		.nios2_instruction_master_readdata               (nios2_instruction_master_readdata),                         //                                          .readdata
		.nios2_instruction_master_readdatavalid          (nios2_instruction_master_readdatavalid),                    //                                          .readdatavalid
		.alarm_select_s1_address                         (mm_interconnect_0_alarm_select_s1_address),                 //                           alarm_select_s1.address
		.alarm_select_s1_write                           (mm_interconnect_0_alarm_select_s1_write),                   //                                          .write
		.alarm_select_s1_readdata                        (mm_interconnect_0_alarm_select_s1_readdata),                //                                          .readdata
		.alarm_select_s1_writedata                       (mm_interconnect_0_alarm_select_s1_writedata),               //                                          .writedata
		.alarm_select_s1_chipselect                      (mm_interconnect_0_alarm_select_s1_chipselect),              //                                          .chipselect
		.epcs_flash_epcs_control_port_address            (mm_interconnect_0_epcs_flash_epcs_control_port_address),    //              epcs_flash_epcs_control_port.address
		.epcs_flash_epcs_control_port_write              (mm_interconnect_0_epcs_flash_epcs_control_port_write),      //                                          .write
		.epcs_flash_epcs_control_port_read               (mm_interconnect_0_epcs_flash_epcs_control_port_read),       //                                          .read
		.epcs_flash_epcs_control_port_readdata           (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                                          .readdata
		.epcs_flash_epcs_control_port_writedata          (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                                          .writedata
		.epcs_flash_epcs_control_port_chipselect         (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                                          .chipselect
		.jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //               jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.laser_fifo_in_csr_address                       (mm_interconnect_0_laser_fifo_in_csr_address),               //                         laser_fifo_in_csr.address
		.laser_fifo_in_csr_write                         (mm_interconnect_0_laser_fifo_in_csr_write),                 //                                          .write
		.laser_fifo_in_csr_read                          (mm_interconnect_0_laser_fifo_in_csr_read),                  //                                          .read
		.laser_fifo_in_csr_readdata                      (mm_interconnect_0_laser_fifo_in_csr_readdata),              //                                          .readdata
		.laser_fifo_in_csr_writedata                     (mm_interconnect_0_laser_fifo_in_csr_writedata),             //                                          .writedata
		.laser_fifo_out_address                          (mm_interconnect_0_laser_fifo_out_address),                  //                            laser_fifo_out.address
		.laser_fifo_out_read                             (mm_interconnect_0_laser_fifo_out_read),                     //                                          .read
		.laser_fifo_out_readdata                         (mm_interconnect_0_laser_fifo_out_readdata),                 //                                          .readdata
		.laser_fifo_out_waitrequest                      (mm_interconnect_0_laser_fifo_out_waitrequest),              //                                          .waitrequest
		.led_timer_s1_address                            (mm_interconnect_0_led_timer_s1_address),                    //                              led_timer_s1.address
		.led_timer_s1_write                              (mm_interconnect_0_led_timer_s1_write),                      //                                          .write
		.led_timer_s1_readdata                           (mm_interconnect_0_led_timer_s1_readdata),                   //                                          .readdata
		.led_timer_s1_writedata                          (mm_interconnect_0_led_timer_s1_writedata),                  //                                          .writedata
		.led_timer_s1_chipselect                         (mm_interconnect_0_led_timer_s1_chipselect),                 //                                          .chipselect
		.nios2_debug_mem_slave_address                   (mm_interconnect_0_nios2_debug_mem_slave_address),           //                     nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write                     (mm_interconnect_0_nios2_debug_mem_slave_write),             //                                          .write
		.nios2_debug_mem_slave_read                      (mm_interconnect_0_nios2_debug_mem_slave_read),              //                                          .read
		.nios2_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_debug_mem_slave_readdata),          //                                          .readdata
		.nios2_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_debug_mem_slave_writedata),         //                                          .writedata
		.nios2_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_debug_mem_slave_byteenable),        //                                          .byteenable
		.nios2_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),       //                                          .waitrequest
		.nios2_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),       //                                          .debugaccess
		.onchip_memory_s1_address                        (mm_interconnect_0_onchip_memory_s1_address),                //                          onchip_memory_s1.address
		.onchip_memory_s1_write                          (mm_interconnect_0_onchip_memory_s1_write),                  //                                          .write
		.onchip_memory_s1_readdata                       (mm_interconnect_0_onchip_memory_s1_readdata),               //                                          .readdata
		.onchip_memory_s1_writedata                      (mm_interconnect_0_onchip_memory_s1_writedata),              //                                          .writedata
		.onchip_memory_s1_byteenable                     (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                          .byteenable
		.onchip_memory_s1_chipselect                     (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                          .chipselect
		.onchip_memory_s1_clken                          (mm_interconnect_0_onchip_memory_s1_clken),                  //                                          .clken
		.power_led_s1_address                            (mm_interconnect_0_power_led_s1_address),                    //                              power_led_s1.address
		.power_led_s1_write                              (mm_interconnect_0_power_led_s1_write),                      //                                          .write
		.power_led_s1_readdata                           (mm_interconnect_0_power_led_s1_readdata),                   //                                          .readdata
		.power_led_s1_writedata                          (mm_interconnect_0_power_led_s1_writedata),                  //                                          .writedata
		.power_led_s1_chipselect                         (mm_interconnect_0_power_led_s1_chipselect),                 //                                          .chipselect
		.protocol_fifo_in_address                        (mm_interconnect_0_protocol_fifo_in_address),                //                          protocol_fifo_in.address
		.protocol_fifo_in_write                          (mm_interconnect_0_protocol_fifo_in_write),                  //                                          .write
		.protocol_fifo_in_writedata                      (mm_interconnect_0_protocol_fifo_in_writedata),              //                                          .writedata
		.protocol_fifo_in_waitrequest                    (mm_interconnect_0_protocol_fifo_in_waitrequest),            //                                          .waitrequest
		.protocol_fifo_in_csr_address                    (mm_interconnect_0_protocol_fifo_in_csr_address),            //                      protocol_fifo_in_csr.address
		.protocol_fifo_in_csr_write                      (mm_interconnect_0_protocol_fifo_in_csr_write),              //                                          .write
		.protocol_fifo_in_csr_read                       (mm_interconnect_0_protocol_fifo_in_csr_read),               //                                          .read
		.protocol_fifo_in_csr_readdata                   (mm_interconnect_0_protocol_fifo_in_csr_readdata),           //                                          .readdata
		.protocol_fifo_in_csr_writedata                  (mm_interconnect_0_protocol_fifo_in_csr_writedata),          //                                          .writedata
		.SCL_s1_address                                  (mm_interconnect_0_scl_s1_address),                          //                                    SCL_s1.address
		.SCL_s1_write                                    (mm_interconnect_0_scl_s1_write),                            //                                          .write
		.SCL_s1_readdata                                 (mm_interconnect_0_scl_s1_readdata),                         //                                          .readdata
		.SCL_s1_writedata                                (mm_interconnect_0_scl_s1_writedata),                        //                                          .writedata
		.SCL_s1_chipselect                               (mm_interconnect_0_scl_s1_chipselect),                       //                                          .chipselect
		.SDA_s1_address                                  (mm_interconnect_0_sda_s1_address),                          //                                    SDA_s1.address
		.SDA_s1_write                                    (mm_interconnect_0_sda_s1_write),                            //                                          .write
		.SDA_s1_readdata                                 (mm_interconnect_0_sda_s1_readdata),                         //                                          .readdata
		.SDA_s1_writedata                                (mm_interconnect_0_sda_s1_writedata),                        //                                          .writedata
		.SDA_s1_chipselect                               (mm_interconnect_0_sda_s1_chipselect),                       //                                          .chipselect
		.spird_fifo_in_csr_address                       (mm_interconnect_0_spird_fifo_in_csr_address),               //                         spird_fifo_in_csr.address
		.spird_fifo_in_csr_write                         (mm_interconnect_0_spird_fifo_in_csr_write),                 //                                          .write
		.spird_fifo_in_csr_read                          (mm_interconnect_0_spird_fifo_in_csr_read),                  //                                          .read
		.spird_fifo_in_csr_readdata                      (mm_interconnect_0_spird_fifo_in_csr_readdata),              //                                          .readdata
		.spird_fifo_in_csr_writedata                     (mm_interconnect_0_spird_fifo_in_csr_writedata),             //                                          .writedata
		.spird_fifo_out_address                          (mm_interconnect_0_spird_fifo_out_address),                  //                            spird_fifo_out.address
		.spird_fifo_out_read                             (mm_interconnect_0_spird_fifo_out_read),                     //                                          .read
		.spird_fifo_out_readdata                         (mm_interconnect_0_spird_fifo_out_readdata),                 //                                          .readdata
		.spird_fifo_out_waitrequest                      (mm_interconnect_0_spird_fifo_out_waitrequest),              //                                          .waitrequest
		.spiwr_fifo_in_address                           (mm_interconnect_0_spiwr_fifo_in_address),                   //                             spiwr_fifo_in.address
		.spiwr_fifo_in_write                             (mm_interconnect_0_spiwr_fifo_in_write),                     //                                          .write
		.spiwr_fifo_in_writedata                         (mm_interconnect_0_spiwr_fifo_in_writedata),                 //                                          .writedata
		.spiwr_fifo_in_waitrequest                       (mm_interconnect_0_spiwr_fifo_in_waitrequest),               //                                          .waitrequest
		.spiwr_fifo_in_csr_address                       (mm_interconnect_0_spiwr_fifo_in_csr_address),               //                         spiwr_fifo_in_csr.address
		.spiwr_fifo_in_csr_write                         (mm_interconnect_0_spiwr_fifo_in_csr_write),                 //                                          .write
		.spiwr_fifo_in_csr_read                          (mm_interconnect_0_spiwr_fifo_in_csr_read),                  //                                          .read
		.spiwr_fifo_in_csr_readdata                      (mm_interconnect_0_spiwr_fifo_in_csr_readdata),              //                                          .readdata
		.spiwr_fifo_in_csr_writedata                     (mm_interconnect_0_spiwr_fifo_in_csr_writedata),             //                                          .writedata
		.status_led_s1_address                           (mm_interconnect_0_status_led_s1_address),                   //                             status_led_s1.address
		.status_led_s1_write                             (mm_interconnect_0_status_led_s1_write),                     //                                          .write
		.status_led_s1_readdata                          (mm_interconnect_0_status_led_s1_readdata),                  //                                          .readdata
		.status_led_s1_writedata                         (mm_interconnect_0_status_led_s1_writedata),                 //                                          .writedata
		.status_led_s1_chipselect                        (mm_interconnect_0_status_led_s1_chipselect),                //                                          .chipselect
		.sysid_control_slave_address                     (mm_interconnect_0_sysid_control_slave_address),             //                       sysid_control_slave.address
		.sysid_control_slave_readdata                    (mm_interconnect_0_sysid_control_slave_readdata),            //                                          .readdata
		.w5500_cs_s1_address                             (mm_interconnect_0_w5500_cs_s1_address),                     //                               w5500_cs_s1.address
		.w5500_cs_s1_write                               (mm_interconnect_0_w5500_cs_s1_write),                       //                                          .write
		.w5500_cs_s1_readdata                            (mm_interconnect_0_w5500_cs_s1_readdata),                    //                                          .readdata
		.w5500_cs_s1_writedata                           (mm_interconnect_0_w5500_cs_s1_writedata),                   //                                          .writedata
		.w5500_cs_s1_chipselect                          (mm_interconnect_0_w5500_cs_s1_chipselect),                  //                                          .chipselect
		.w5500_int_s1_address                            (mm_interconnect_0_w5500_int_s1_address),                    //                              w5500_int_s1.address
		.w5500_int_s1_write                              (mm_interconnect_0_w5500_int_s1_write),                      //                                          .write
		.w5500_int_s1_readdata                           (mm_interconnect_0_w5500_int_s1_readdata),                   //                                          .readdata
		.w5500_int_s1_writedata                          (mm_interconnect_0_w5500_int_s1_writedata),                  //                                          .writedata
		.w5500_int_s1_chipselect                         (mm_interconnect_0_w5500_int_s1_chipselect),                 //                                          .chipselect
		.w5500_rst_s1_address                            (mm_interconnect_0_w5500_rst_s1_address),                    //                              w5500_rst_s1.address
		.w5500_rst_s1_write                              (mm_interconnect_0_w5500_rst_s1_write),                      //                                          .write
		.w5500_rst_s1_readdata                           (mm_interconnect_0_w5500_rst_s1_readdata),                   //                                          .readdata
		.w5500_rst_s1_writedata                          (mm_interconnect_0_w5500_rst_s1_writedata),                  //                                          .writedata
		.w5500_rst_s1_chipselect                         (mm_interconnect_0_w5500_rst_s1_chipselect)                  //                                          .chipselect
	);

	kernel_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
